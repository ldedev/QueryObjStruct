module contracts

pub interface IToken {
mut:
	value string
	typ TypeToken
}
