module contracts

pub enum TypeToken {
	undefined
	key
	object
	object_root
	array_all_index
	array_index
	function
}
