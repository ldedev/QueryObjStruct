module contracts
pub interface IArgument {
mut:
	name string
	typ TypeArgument
}
