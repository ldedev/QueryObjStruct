module contracts

pub enum TypeArgument {
	literal
	key
}
