module entities

import contracts { TypeArgument }

pub struct Argument {
pub mut:
	name string
	typ TypeArgument
}
